`timescale 1ns/10ps
module LEDDC( DCK, DAI, DEN, GCK, Vsync, mode, rst, OUT);
input           DCK;
input           DAI;
input           DEN;
input           GCK;
input           Vsync;
input           mode;
input           rst;
output [15:0]   OUT;

// ------------------------------------------------------------
// parameter & genvar
// ------------------------------------------------------------
parameter IDLE     = 5'd17;
parameter CNT_15   = 5'd15;
parameter CNT_14   = 5'd14;
parameter CNT_13   = 5'd13;
parameter CNT_12   = 5'd12;
parameter CNT_11   = 5'd11;
parameter CNT_10   = 5'd10;
parameter CNT_9    = 5'd9;
parameter CNT_8    = 5'd8;
parameter CNT_7    = 5'd7;
parameter CNT_6    = 5'd6;
parameter CNT_5    = 5'd5;
parameter CNT_4    = 5'd4;
parameter CNT_3    = 5'd3;   
parameter CNT_2    = 5'd2;
parameter CNT_1    = 5'd1;
parameter CNT_0    = 5'd0;
parameter CNT_LAST = 5'd16;


genvar i, j;



// ------------------------------------------------------------
// regs & wire
// ------------------------------------------------------------
reg  [15:0] cnt_pwm;
wire [16:0] cnt_pwm_w;
reg  [15:0] pxl_current[15:0], pxl_nxt[15:0];
reg  pwm_sel;

reg [4:0]  cs;
reg cnt_round;


// ------------------------------------------------------------
// design
// ------------------------------------------------------------


always @(posedge GCK or posedge rst) begin
	if (rst) cs <= IDLE;
	else begin
		case (cs)
			IDLE :  cs <= (Vsync) ? ((mode) ? CNT_14 : CNT_15) : IDLE;
			CNT_15: cs <= (pwm_sel) ? CNT_14   : CNT_15;
			CNT_14: cs <= (pwm_sel) ? CNT_13   : CNT_14; 
			CNT_13: cs <= (pwm_sel) ? CNT_12   : CNT_13;
			CNT_12: cs <= (pwm_sel) ? CNT_11   : CNT_12;
			CNT_11: cs <= (pwm_sel) ? CNT_10   : CNT_11;
			CNT_10: cs <= (pwm_sel) ? CNT_9    : CNT_10;
			CNT_9:  cs <= (pwm_sel) ? CNT_8    : CNT_9;
			CNT_8:  cs <= (pwm_sel) ? CNT_7    : CNT_8;
			CNT_7:  cs <= (pwm_sel) ? CNT_6    : CNT_7;
			CNT_6:  cs <= (pwm_sel) ? CNT_5    : CNT_6;
			CNT_5:  cs <= (pwm_sel) ? CNT_4    : CNT_5;
			CNT_4:  cs <= (pwm_sel) ? CNT_3    : CNT_4;
			CNT_3:  cs <= (pwm_sel) ? CNT_2    : CNT_3;
			CNT_2:  cs <= (pwm_sel) ? CNT_1    : CNT_2;
			CNT_1:  cs <= (pwm_sel) ? CNT_0    : CNT_1;
			CNT_0:  cs <= (pwm_sel) ? CNT_LAST : CNT_0;
			CNT_LAST: cs <= IDLE;
			default:  cs <= IDLE;
		endcase
	end
end


always @(posedge GCK or posedge rst) begin
	if (rst) cnt_pwm <= 16'd0;
	else	 cnt_pwm <= (pwm_sel) ? 16'd0 : cnt_pwm_w[15:0];
end

assign cnt_pwm_w = cnt_pwm + 16'd1;
always @(*) begin
	case (cs)
		CNT_15: pwm_sel <= (cnt_pwm_w[16]);
		CNT_14: pwm_sel <= (cnt_pwm_w[15]); 
		CNT_13: pwm_sel <= (cnt_pwm_w[14]);
		CNT_12: pwm_sel <= (cnt_pwm_w[13]);
		CNT_11: pwm_sel <= (cnt_pwm_w[12]);
		CNT_10: pwm_sel <= (cnt_pwm_w[11]);
		CNT_9:  pwm_sel <= (cnt_pwm_w[10]);
		CNT_8:  pwm_sel <= (cnt_pwm_w[9]);
		CNT_7:  pwm_sel <= (cnt_pwm_w[8]);
		CNT_6:  pwm_sel <= (cnt_pwm_w[7]);
		CNT_5:  pwm_sel <= (cnt_pwm_w[6]);
		CNT_4:  pwm_sel <= (cnt_pwm_w[5]);
		CNT_3:  pwm_sel <= (cnt_pwm_w[4]);
		CNT_2:  pwm_sel <= (cnt_pwm_w[3]);
		CNT_1:  pwm_sel <= (cnt_pwm_w[2]);
		CNT_0:  pwm_sel <= (cnt_pwm_w[1]);
		default:  pwm_sel <= 1'b0;
	endcase
end


always @(posedge GCK or posedge rst) begin
	if (rst) cnt_round <= 1'b0;
	else 	 cnt_round <= (cs == CNT_LAST && mode) ? !cnt_round : cnt_round;
end

generate 
for (i = 0; i < 16; i = i + 1) begin
	for (j = 0; j < 16; j = j + 1) begin
		if (j == 0) begin
			always @(posedge GCK or posedge rst) begin
				if (rst) 	     pxl_current[i][j] <= 1'b0;
				else if (!Vsync) pxl_current[i][j] <= (round || !mode) ? 1'b0 : pxl_nxt[i][0];
				else 	 	     pxl_current[i][j] <= pxl_current[i][j];
			end
		end
		else begin
			always @(posedge GCK or posedge rst) begin
				if (rst) 			 			pxl_current <= 16'd0;
				else if (!Vsync)     			pxl_current[i][j] <= pxl_nxt[i][j];
 				else if (cs != IDLE && pwm_sel) pxl_current[i][j] <= pxl_current[i][j - 1];
				else 	 			 			pxl_current[i][j] <= pxl_current[i][j];
			end
		end
	end

end
endgenerate


generate 
for (i = 0; i < 16; i = i + 1) begin
	always @(posedge GCK or posedge rst) begin
		if (rst) OUT[i] <= 1'b0;
		else  	 OUT[i] <= (Vsync) ? pxl_current[i][15] : 1'b0;
	end
end
endgenerate

endmodule
